module ALU(mode, a, b, o);
    assign [3:0] mode;
    input [3:0]a,b ;
    output [3:0]o;

